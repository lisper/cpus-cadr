/*
 * $Id$
 */

module part_74S241(AENB_N, BENB,
		   Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7);

  input AENB_N, BENB;
  output Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7;

endmodule

/*
 * $Id$
 */

module part_74S157 ( A1, B1, A2, B2, A3, B3, B4, A4, 
		     Y1, Y2, Y3, Y4,
		     SEL, ENB_N );
  input A1, B1, A2, B2, A3, B3, B4, A4;
  output Y1, Y2, Y3, Y4;
  input SEL, ENB_N;

endmodule

/*
 * $Id$
 */

module part_9S42_1 ( G1A1, G1B1, G2A1, G2B1, G2C1, G2D1, 
		     G1A2, G1B2, G2A2, G2B2, G2C2, G2D2,
		     OUT1, OUT2 );
  input G1A1, G1B1, G2A1, G2B1, G2C1, G2D1;
  input G1A2, G1B2, G2A2, G2B2, G2C2, G2D2;
  output OUT1, OUT2;

  assign OUT1 = (G1A1 & G1B1) | (G2A1 & G2B1 & G2C1 & G2D1);
  assign OUT2 = (G1A2 & G1B2) | (G2A2 & G2B2 & G2C2 & G2D2);

endmodule

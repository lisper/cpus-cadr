/*
 * $Id$
 */

module part_TD50 ( INPUT, O_10ns, O_20ns, O_30ns, O_40ns, O_50ns );
  input INPUT;
  output O_10ns, O_20ns, O_30ns, O_40ns, O_50ns;

endmodule

/*
 * $Id$
 */

module part_74LS244(D0, D1, D2, D3, D4, D5, D6, D7,
		    Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7,
		EN1_N, EN2_N);
  input D0, D1, D2, D3, D4, D5, D6, D7;
  output Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7;
  input EN1_N, EN2_N;

endmodule

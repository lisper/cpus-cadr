/*
 * $Id$
 */

module part_TIL309 (I1, I2, I4, I8, DP, LDP, LATCH, BLANK_N, TEST_N,
	L1, L2, L4, L8);

  input I1, I2, I4, I8, DP, LDP, LATCH, BLANK_N, TEST_N;
  output L1, L2, L4, L8;

endmodule

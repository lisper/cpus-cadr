/*
 * $Id$
 */

module part_2147 (A0,A1,A2,A3,A4,A5,A6,A7,A8,A9,A10,A11, CE_N, WE_N, DI, DO);

  input A0,A1,A2,A3,A4,A5,A6,A7,A8,A9,A10,A11;
  input CE_N, WE_N, DI;
  output DO;

endmodule

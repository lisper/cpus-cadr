/*
 * $Id$
 */

module part_TD100 ( INPUT, O_20ns, O_40ns, O_60ns, O_80ns, O_100ns );
  input INPUT;
  output O_20ns, O_40ns, O_60ns, O_80ns, O_100ns;

endmodule

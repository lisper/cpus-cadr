/*
 * $Id$
 */

module part_74S258 (A0, A1, B0, B1, C0, C1, D0, D1,
		SEL, ENB_N, AY, BY, CY, DY);

  input A0, A1, B0, B1, C0, C1, D0, D1;
  input SEL, ENB_N;
  output AY, BY, CY, DY;

endmodule


module part_16DUMMY ();

endmodule

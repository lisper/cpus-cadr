/*
 * $Id$
 */

module part_SIP330_470_8 (R2, R3, R4, R5, R6, R7);
  output R2, R3, R4, R5, R6, R7;

  pullup p2(R2);
  pullup p3(R3);
  pullup p4(R4);
  pullup p5(R5);
  pullup p6(R6);
  pullup p7(R7);

endmodule

module part_SIP220_330_8(R2, R3, R4, R5, R6, R7);
  output R2, R3, R4, R5, R6, R7;

  pullup p2(R2);
  pullup p3(R3);
  pullup p4(R4);
  pullup p5(R5);
  pullup p6(R6);
  pullup p7(R7);

endmodule
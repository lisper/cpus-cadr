/*
 * $Id$
 */

module part_74S174 (D1, Q1, D2, Q2, D3, Q3, D4, Q4, D5, Q5, D6, Q6,
	CLR_N, CLK);

  input D1, D2, D3, D4, D5, D6;
  input CLR_N, CLK;
  output Q1, Q2, Q3, Q4, Q5, Q6;

endmodule

/*
 * $Id$
 */

module part_74S175 (D0, Q0, Q0_N, D1, Q1, Q1_N, D2, Q2, Q2_N, D3, Q3, Q3_N,
	CLR_N, CLK);

  input D0, D1, D2, D3;
  input CLR_N, CLK;
  output Q0, Q0_N, Q1, Q1_N, Q2, Q2_N, Q3, Q3_N;

endmodule

/*
 * $Id$
 */

module part_93S48(I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, PE, PO);

  input I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11;
  output PE, PO;

endmodule

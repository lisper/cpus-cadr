/*
 * $Id$
 */

module part_25S10 (I3, I2, I1, I0, I_1, I_2, I_3,
	SEL0, SEL1, CE_N,
	O0, O1, O2, O3);

  input I3, I2, I1, I0, I_1, I_2, I_3;
  input SEL0, SEL1, CE_N;
  output O0, O1, O2, O3;

endmodule

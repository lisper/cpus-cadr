/*
 * $Id$
 */

module part_74S153 ( G1D0, G1D1, G1D2, G1D3,
		     G2D0, G2D1, G2D2, G2D3,
		     G1Q, G2Q,
		     SEL0, SEL1, ENB1_N, ENB2_N);

  input G1D0, G1D1, G1D2, G1D3;
  input G2D0, G2D1, G2D2, G2D3;

  input SEL0, SEL1, ENB1_N, ENB2_N;
  output G1Q, G2Q;

endmodule

/*
 * $Id$
 */

module part_82S21 (I0, I1, A0, A1, A2, A3, A4,
		WE0_N, WE1_N, LATCH_N, WCLK_N, CE,
		D0, D1);

  input I0, I1, A0, A1, A2, A3, A4;
  input WE0_N, WE1_N, LATCH_N, WCLK_N, CE;
  output D0, D1;

endmodule

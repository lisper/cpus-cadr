/*
 * $Id$
 */

module part_RES20(R2, R3, R4, R5, R6, R7, R8, R9, R10,
		  R11, R12, R13, R14, R15, R16, R17, R18, R19);
  output R2, R3, R4, R5, R6, R7, R8, R9, R10;
  output R11, R12, R13, R14, R15, R16, R17, R18, R19;

/*  assign R2 = pullup; */

endmodule

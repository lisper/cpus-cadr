/*
 * $Id$
 */

module part_TD250 ( INPUT, O_50ns, O_100ns, O_150ns, O_200ns, O_250ns );
  input INPUT;
  output O_50ns, O_100ns, O_150ns, O_200ns, O_250ns;

endmodule

/*
 * $Id$
 */

module part_SIP330_470_8 (R2, R3, R4, R5, R6, R7);
  input R2, R3, R4, R5, R6, R7;

endmodule

module part_SIP220_330_8(R2, R3, R4, R5, R6, R7);
  input R2, R3, R4, R5, R6, R7;
endmodule

module part_16DUMMY (dummy);
  input dummy;

endmodule

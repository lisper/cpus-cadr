/*
 * $Id$
 */

module part_74S74 ( G1R_N, G1D, G1CLK, G1S_N, G2S_N, G2CLK, G2D, G2R_N,
	G1Q, G1Q_N, G2Q_N, G2Q);

  input G1R_N, G1D, G1CLK, G1S_N;
  input G2S_N, G2CLK, G2D, G2R_N;
  output G1Q, G1Q_N, G2Q_N, G2Q;

endmodule

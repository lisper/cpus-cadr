/*
 * $Id$
 */

module part_74S280 (I0, I1, I2, I3, I4, I5, I6, I7, I8,
	EVEN, ODD);

  input I0, I1, I2, I3, I4, I5, I6, I7, I8;
  output EVEN, ODD;

endmodule

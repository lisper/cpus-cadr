/*
 * $Id$
 */

module part_74S169 (I0, I1, I2, I3,
	O3, O2, O1, O0,
	CO_N, ENB_T_N, ENB_P_N, LOAD_N, UP_DN, CLK);

  input I0, I1, I2, I3;
  output O3, O2, O1, O0;
  input CO_N, ENB_T_N, ENB_P_N, LOAD_N, UP_DN, CLK;

endmodule

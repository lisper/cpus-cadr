/*
 * $Id$
 */

module part_TD25 ( INPUT, O_5ns, O_10ns, O_15ns, O_20ns, O_25ns );
  input INPUT;
  output O_5ns, O_10ns, O_15ns, O_20ns, O_25ns;

endmodule

/*
 * $Id$
 */

module part_74S194 (I0, I1, I2, I3,
	Q3, Q2, Q1, Q0,
	CLR_N, SIL, SIR, S0, S1, CLK);

  input I0, I1, I2, I3;
  output Q3, Q2, Q1, Q0;
  input CLR_N, SIL, SIR, S0, S1, CLK;

endmodule

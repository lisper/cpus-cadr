/*
 * $Id$
 */

module part_74S139( A1, B1, G1,
	A2, B2, G2,
	G1Y0, G1Y1, G1Y2, G1Y3, G2Y0, G2Y1, G2Y2, G2Y3);

  input A1, B1, G1;
  input A2, B2, G2;
  output G1Y0, G1Y1, G1Y2, G1Y3, G2Y0, G2Y1, G2Y2, G2Y3;

endmodule
